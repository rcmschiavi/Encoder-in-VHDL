

entity gerenciador is
	port(
		dir: in std_logic;
		cont: in std_logic_vector(6 downto 0);
		dado: out std_logic_vector(7 downto 0);
	);
end gerenciador;

architecture gerenciamento of gerenciador is


	begin
	
		
	
end gerenciamento	