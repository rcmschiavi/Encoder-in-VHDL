

entity gerenciador is
	port(
		dir: in
	);
end gerenciador;

architecture gerenciamento of gerenciador is


	begin
	
		
	
end gerenciamento	